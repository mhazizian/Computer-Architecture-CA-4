`include "defines.sv"

module PR_1_IF_ID(clk, rst, PR1_PC_plus1, PR1_instruction_in, PC_plus1, instruction);
	input clk, rst;
	input [`INSTRUCTION_LEN - 1:0] PR1_instruction_in;
	input [`ADDRESS_LEN - 1:0] PR1_PC_plus1;

	output logic [`INSTRUCTION_LEN - 1:0] PR1_Instruction;
	output logic [`ADDRESS_LEN - 1:0] PC_plus1;

	always@(posedge clk, posedge rst) begin
		if(rst) begin
			PC_plus1 <= 0;
			instruction <= 0;
		end
		else begin
			PC_plus1 <= PR1_PC_plus1;
			instruction <= PR1_instruction_in;
		end
	end
endmodule // PR_1_IF_ID